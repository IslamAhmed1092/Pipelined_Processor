library ieee; 
use ieee.std_logic_1164.all; 
USE IEEE.numeric_std.all;

entity control_store is 
port (out_data: out std_logic_vector(31 downto 0); 
    address: In std_logic_vector(8 downto 0));
end control_store; 

architecture control_store_arc of control_store is 
type control_store_type is array (0 to 511) of std_logic_vector(31 downto 0); 

SIGNAL control_store : control_store_type := (
    -- F0   Next instruction
    -- F1   No,PC,MDR,Z,Rs,Rd,S,D,T,Address     Out        
    -- F2   No,PC,IR,Z,Rs,Rd                    IN 
    -- F3   No,MAR,MDR,TEMP                     IN
    -- F4   No,Y,S,D                            IN
    -- F5   MOV,ADD,ADC,SUB,SBC,AND,OR,XOR,CMP,INC,DEC,CLR,INV,LSR,ROR,ASR,LSL,ROL
    -- F6   No,READ,WRITE,CLOCK_ENABLE
    -- F7   No,WMFC
    -- F8   No,ORdst,ORindsrc,ORinddst,ORresult,ORoperations
    -- F9   No,PLAout
    
    --------------------------------------START------------------------------------------------
    --      "F0"     "F1"    "F2"    "F3"   "F4"     "F5"   "F6"   "F7"  "F8"    "F9"
    0   => o"001" & "0001" & "011" & "01" & "01" & "01001" & "01" & "0" & "000" & "0",
    1   => o"002" & "0011" & "001" & "00" & "00" & "00000" & "00" & "1" & "000" & "0",
    2   => o"003" & "0010" & "010" & "00" & "00" & "00000" & "00" & "0" & "000" & "0",
    3   => o"000" & "0000" & "000" & "00" & "00" & "00000" & "00" & "0" & "000" & "1",

    
   
    -----------------------------------2&1 operands--------------------------------------------
    
    ----------------------------------fetcing source-------------------------------------------
    272 => o"470" & "0100" & "000" & "00" & "10" & "00000" & "00" & "0" & "001" & "0",
    
    280 => o"466" & "0100" & "000" & "01" & "00" & "00000" & "01" & "1" & "000" & "0",
    
    288 => o"441" & "0100" & "011" & "01" & "01" & "01001" & "01" & "0" & "000" & "0",
    289 => o"465" & "0011" & "100" & "00" & "00" & "00000" & "01" & "1" & "010" & "0",
 
    296 => o"451" & "0100" & "011" & "00" & "01" & "01010" & "00" & "0" & "000" & "0",
    297 => o"465" & "0011" & "100" & "01" & "00" & "00000" & "01" & "1" & "010" & "0",

    304 => o"461" & "0001" & "011" & "01" & "01" & "01001" & "01" & "0" & "000" & "0",
    305 => o"462" & "0011" & "001" & "00" & "00" & "00000" & "00" & "1" & "000" & "0",
    306 => o"463" & "0010" & "000" & "00" & "01" & "00000" & "00" & "0" & "000" & "0",
    307 => o"464" & "0100" & "011" & "00" & "00" & "00001" & "00" & "0" & "000" & "0",
    308 => o"465" & "0011" & "000" & "01" & "00" & "00000" & "01" & "1" & "010" & "0",


    309 => o"466" & "0010" & "000" & "01" & "00" & "00000" & "01" & "1" & "000" & "0",
    310 => o"470" & "0010" & "000" & "00" & "10" & "00000" & "00" & "0" & "001" & "0",



    ----------------------------------fetcing destination-------------------------------------------

    312 => o"537" & "0101" & "000" & "00" & "01" & "00000" & "00" & "0" & "101" & "0",
    
    320 => o"536" & "0101" & "000" & "01" & "00" & "00000" & "01" & "1" & "000" & "0",
    
    328 => o"511" & "0101" & "011" & "01" & "01" & "01001" & "01" & "0" & "000" & "0",
    329 => o"535" & "0011" & "101" & "00" & "00" & "00000" & "01" & "1" & "011" & "0",
 
    336 => o"521" & "0101" & "011" & "00" & "01" & "01010" & "00" & "0" & "000" & "0",
    337 => o"535" & "0011" & "101" & "01" & "00" & "00000" & "01" & "1" & "011" & "0",

    344 => o"531" & "0001" & "011" & "01" & "01" & "01001" & "01" & "0" & "000" & "0",
    345 => o"532" & "0011" & "001" & "00" & "00" & "00000" & "00" & "1" & "000" & "0",
    346 => o"533" & "0010" & "000" & "00" & "01" & "00000" & "00" & "0" & "000" & "0",
    347 => o"534" & "0101" & "011" & "00" & "01" & "00001" & "00" & "0" & "000" & "0",
    348 => o"535" & "0011" & "000" & "01" & "00" & "00000" & "01" & "1" & "011" & "0",

    349 => o"536" & "0010" & "000" & "01" & "00" & "00000" & "01" & "1" & "000" & "0",
    350 => o"537" & "0010" & "000" & "00" & "01" & "00000" & "00" & "0" & "101" & "0",

    351 => o"561" & "1000" & "011" & "00" & "00" & "00000" & "00" & "0" & "100" & "0",
    352 => o"561" & "1000" & "011" & "00" & "00" & "00001" & "00" & "0" & "100" & "0",
    353 => o"561" & "1000" & "011" & "00" & "00" & "00010" & "00" & "0" & "100" & "0",
    354 => o"561" & "1000" & "011" & "00" & "00" & "00011" & "00" & "0" & "100" & "0",
    355 => o"561" & "1000" & "011" & "00" & "00" & "00100" & "00" & "0" & "100" & "0",
    356 => o"561" & "1000" & "011" & "00" & "00" & "00101" & "00" & "0" & "100" & "0",
    357 => o"561" & "1000" & "011" & "00" & "00" & "00110" & "00" & "0" & "100" & "0",
    358 => o"561" & "1000" & "011" & "00" & "00" & "00111" & "00" & "0" & "100" & "0",
    359 => o"000" & "1000" & "011" & "00" & "00" & "01000" & "00" & "0" & "100" & "0",
    360 => o"561" & "1000" & "011" & "00" & "00" & "01001" & "00" & "0" & "100" & "0",
    361 => o"561" & "1000" & "011" & "00" & "00" & "01010" & "00" & "0" & "100" & "0",
    362 => o"561" & "1000" & "011" & "00" & "00" & "01011" & "00" & "0" & "100" & "0",
    363 => o"561" & "1000" & "011" & "00" & "00" & "01100" & "00" & "0" & "100" & "0",
    364 => o"561" & "1000" & "011" & "00" & "00" & "01101" & "00" & "0" & "100" & "0",
    365 => o"561" & "1000" & "011" & "00" & "00" & "01110" & "00" & "0" & "100" & "0",
    366 => o"561" & "1000" & "011" & "00" & "00" & "01111" & "00" & "0" & "100" & "0",
    367 => o"561" & "1000" & "011" & "00" & "00" & "10000" & "00" & "0" & "100" & "0",
    368 => o"561" & "1000" & "011" & "00" & "00" & "10001" & "00" & "0" & "100" & "0",


    369 => o"000" & "0011" & "000" & "10" & "00" & "00000" & "10" & "0" & "000" & "0",
    370 => o"000" & "0011" & "101" & "00" & "00" & "00000" & "00" & "0" & "000" & "0",




    -------------------------------------branching---------------------------------------------
    184 => o"271" & "0001" & "000" & "00" & "01" & "00000" & "00" & "0" & "000" & "0",
    185 => o"272" & "1011" & "011" & "00" & "00" & "00001" & "00" & "0" & "000" & "0",
    186 => o"000" & "0011" & "001" & "00" & "00" & "00000" & "00" & "0" & "000" & "0",


    -------------------------------------No Operand--------------------------------------------
    96 => o"141" & "0001" & "011" & "00" & "01" & "01001" & "00" & "0" & "000" & "0",
    97 => o"000" & "0011" & "001" & "00" & "00" & "00000" & "00" & "0" & "000" & "0",
    98 => o"000" & "0000" & "000" & "00" & "00" & "00000" & "11" & "0" & "000" & "0",
    


    
    others => x"00000000"
);

begin
    out_data <= control_store(to_integer(unsigned(address)));
end control_store_arc; 
    